`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// vga_driver.v -- basic video driver
//
// Author:  W. Freund, UTFSM, Valparaiso, Chile
//          (based on vga_main.vhd from Barron Barnett, Digilent, Inc.) 
//          03/05/06, 14/06/12
//Modifier: Mauricio Solis
//				28/05/2014
//Modifier: Mauricio Solis
//				09/06/2017
////////////////////////////////////////////////////////////////////////////////
//http://tinyvga.com/vga-timing/800x600@72Hz

module driver_vga_1024x768(
		input clk_vga,
        input rst,                    
		output hs, vs,
		output [10:0]hc_visible,
        output [10:0]vc_visible
        ); 
    
        //1024x768 @60Hz XGA
        localparam hpixels = 11'd1344;  // --Value of pixels in a horizontal line
        localparam vlines  = 11'd806
        ;  // --Number of horizontal lines in the display
    
        localparam hfp  = 11'd24;      // --Horizontal front porch
        localparam hsc  = 11'd136;      // --Horizontal sync
        localparam hbp  = 11'd160;      // --Horizontal back porch
        
        localparam vfp  = 11'd3;       // --Vertical front porch
        localparam vsc  = 11'd6;       // --Vertical sync
        localparam vbp  = 11'd29;      // --Vertical back porch
        
        
        logic [10:0] hc, hc_next, vc, vc_next;             // --These are the Horizontal and Vertical counters    
        
        assign hc_visible = ((hc < (hpixels - hfp+1)) && (hc > (hsc + hbp)))?(hc -(hsc + hbp)):10'd0;
        assign vc_visible = ((vc < (vlines - vfp+1)) && (vc > (vsc + vbp)))?(vc - (vsc + vbp)):10'd0;
        
        
        // --Runs the horizontal counter
    
        always_comb
            if(hc == hpixels)                // --If the counter has reached the end of pixel count
                hc_next = 11'd0;            // --reset the counter
            else
                hc_next = hc + 11'd1;        // --Increment the horizontal counter
    
        
        // --Runs the vertical counter
        always_comb
            if(hc == 11'd0)
                if(vc == vlines)
                    vc_next = 11'd0;
                else
                    vc_next = vc + 11'd1;
            else
                vc_next = vc;
        
        always_ff@(posedge clk_vga)
            if (rst)
                {hc, vc} <= 'd0;
            else
                {hc, vc} <= {hc_next, vc_next};
            
        assign hs = (hc < hsc) ? 1'b0 : 1'b1;   // --Horizontal Sync Pulse
        assign vs = (vc < vsc) ? 1'b0 : 1'b1;   // --Vertical Sync Pulse
        
    endmodule